`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/06/28 15:47:02
// Design Name: 
// Module Name: Instr_Decoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Instr_dec(
    input [31:0] instr_code,
    output reg [31:0] code
    );
    wire [11:0] t;
    assign t = {instr_code[31:26],instr_code[5:0]};
    always @ (*)
    begin
        casez(t)
            12'b000000100000 :code = 32'b00000000000000000000000000000001;    //ADD
            12'b000000100001 :code = 32'b00000000000000000000000000000010;    //ADDU
            12'b000000100010 :code = 32'b00000000000000000000000000000100;    //SUB
            12'b000000100011 :code = 32'b00000000000000000000000000001000;    //SUBU
            12'b000000100100 :code = 32'b00000000000000000000000000010000;    //AND
            12'b000000100101 :code = 32'b00000000000000000000000000100000;    //OR
            12'b000000100110 :code = 32'b00000000000000000000000001000000;    //XOR
            12'b000000100111 :code = 32'b00000000000000000000000010000000;    //NOR
            12'b000000101010 :code = 32'b00000000000000000000000100000000;    //SLT
            12'b000000101011 :code = 32'b00000000000000000000001000000000;    //SLTU
            12'b000000000000 :code = 32'b00000000000000000000010000000000;    //SLL
            12'b000000000010 :code = 32'b00000000000000000000100000000000;    //SRL
            12'b000000000011 :code = 32'b00000000000000000001000000000000;    //SRA
            12'b000000000100 :code = 32'b00000000000000000010000000000000;    //SLLV
            12'b000000000110 :code = 32'b00000000000000000100000000000000;    //SRLV
            12'b000000000111 :code = 32'b00000000000000001000000000000000;    //SRAV
            12'b000000001000 :code = 32'b00000000000000010000000000000000;    //JR
            12'b001000?????? :code = 32'b00000000000000100000000000000000;    //ADDI
            12'b001001?????? :code = 32'b00000000000001000000000000000000;    //ADDIU
            12'b001100?????? :code = 32'b00000000000010000000000000000000;    //ANDI
            12'b001101?????? :code = 32'b00000000000100000000000000000000;    //ORI
            12'b001110?????? :code = 32'b00000000001000000000000000000000;    //XORI
            12'b100011?????? :code = 32'b00000000010000000000000000000000;    //LW
            12'b101011?????? :code = 32'b00000000100000000000000000000000;    //SW
            12'b000100?????? :code = 32'b00000001000000000000000000000000;    //BEQ
            12'b000101?????? :code = 32'b00000010000000000000000000000000;    //BNE
            12'b001010?????? :code = 32'b00000100000000000000000000000000;    //SLTI
            12'b001011?????? :code = 32'b00001000000000000000000000000000;    //SLTIU
            12'b001111?????? :code = 32'b00010000000000000000000000000000;    //LUI
            12'b000010?????? :code = 32'b00100000000000000000000000000000;    //J
            12'b000011?????? :code = 32'b01000000000000000000000000000000;    //JAL
            default:          code = 32'bx;
        endcase
    end
    
endmodule
